`ifndef TB_ENV_PKG_SV
`define TB_ENV_PKG_SV
package tb_env_pkg;
  import  uvm_pkg::*;
  import  tue_pkg::*;
  import  tvip_common_pkg::*;
  import  tvip_apb_pkg::*;
  import  sample_0_ral_pkg::*;
  import  sample_1_ral_pkg::*;

  `include  "uvm_macros.svh"
  `include  "tue_macros.svh"

  `include  "tb_env_configuration.svh"
  `include  "tb_env_ral_model.svh"
  `include  "tb_env_ral.svh"
  `include  "tb_env.svh"
endpackage
`endif
