`ifndef TB_ENV_RAL_MODEL_SVH
`define TB_ENV_RAL_MODEL_SVH
class tb_env_ral_model extends sample_0_block_model #(sample_1_block_model);
  `tue_object_default_constructor(tb_env_ral_model)
  `uvm_object_utils(tb_env_ral_model)
endclass
`endif
